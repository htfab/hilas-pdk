VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_fgvaractorcapacitor02
  CLASS BLOCK ;
  FOREIGN sky130_hilas_fgvaractorcapacitor02 ;
  ORIGIN 10.050 3.800 ;
  SIZE 2.720 BY 1.690 ;
  OBS
      LAYER nwell ;
        RECT -10.050 -2.150 -7.340 -2.110 ;
        RECT -10.050 -3.800 -7.330 -2.150 ;
      LAYER li1 ;
        RECT -9.750 -3.280 -9.520 -2.590 ;
      LAYER mcon ;
        RECT -9.720 -2.800 -9.550 -2.630 ;
        RECT -9.720 -3.250 -9.550 -3.080 ;
      LAYER met1 ;
        RECT -9.770 -3.330 -9.510 -2.540 ;
  END
END sky130_hilas_fgvaractorcapacitor02
END LIBRARY

