magic
tech sky130A
timestamp 1634057717
<< checkpaint >>
rect 821 1716 2254 1720
rect 702 1547 2254 1716
rect 702 1362 2654 1547
rect 410 101 2654 1362
rect 410 -189 2254 101
rect 410 -194 2185 -189
rect 410 -630 1926 -194
<< error_s >>
rect 818 657 868 663
rect 890 657 940 663
rect 818 615 868 621
rect 890 615 940 621
rect 818 588 868 594
rect 818 546 868 552
rect 818 503 868 509
rect 818 461 868 467
rect 818 434 868 440
rect 890 434 940 440
rect 818 392 868 398
rect 890 392 940 398
rect 818 333 868 339
rect 890 333 940 339
rect 818 291 868 297
rect 890 291 940 297
rect 818 264 868 270
rect 818 222 868 228
rect 818 180 868 186
rect 818 138 868 144
rect 818 111 868 117
rect 890 111 940 117
rect 818 69 868 75
rect 890 69 940 75
<< nwell >>
rect 0 557 7 575
rect 57 522 116 533
rect 431 516 542 539
rect 895 373 930 374
rect 895 357 912 373
rect 929 357 930 373
rect 57 194 116 213
rect 431 192 542 219
<< psubdiff >>
rect 278 527 304 550
rect 278 510 282 527
rect 299 510 304 527
rect 670 526 697 552
rect 278 484 304 510
rect 670 509 676 526
rect 693 509 697 526
rect 670 486 697 509
rect 279 415 304 442
rect 279 398 283 415
rect 300 398 304 415
rect 279 381 304 398
rect 279 364 283 381
rect 300 364 304 381
rect 279 347 304 364
rect 279 330 283 347
rect 300 330 304 347
rect 279 302 304 330
rect 672 401 697 428
rect 672 384 676 401
rect 693 384 697 401
rect 672 367 697 384
rect 672 350 676 367
rect 693 350 697 367
rect 672 333 697 350
rect 672 316 676 333
rect 693 316 697 333
rect 672 303 697 316
<< mvnsubdiff >>
rect 57 522 116 533
rect 431 516 542 539
rect 57 194 116 213
rect 431 192 542 219
<< psubdiffcont >>
rect 282 510 299 527
rect 676 509 693 526
rect 283 398 300 415
rect 283 364 300 381
rect 283 330 300 347
rect 676 384 693 401
rect 676 350 693 367
rect 676 316 693 333
<< poly >>
rect 583 596 751 613
rect 156 559 393 583
rect 156 450 391 474
rect 582 442 751 459
rect 912 373 930 374
rect 928 357 930 373
rect 156 270 393 294
rect 640 289 660 295
rect 583 272 751 289
rect 158 120 391 144
rect 583 120 752 136
<< polycont >>
rect 895 357 912 374
<< locali >>
rect 282 527 299 529
rect 676 526 693 528
rect 283 415 300 423
rect 283 381 300 383
rect 283 322 300 330
rect 676 401 693 409
rect 676 367 693 369
rect 886 357 895 374
rect 676 308 693 316
<< viali >>
rect 282 529 299 546
rect 282 493 299 510
rect 676 528 693 545
rect 676 492 693 509
rect 283 398 300 400
rect 283 383 300 398
rect 283 347 300 364
rect 676 384 693 386
rect 676 369 693 384
rect 912 357 930 374
rect 676 333 693 350
<< metal1 >>
rect 35 41 75 691
rect 279 550 303 691
rect 440 658 478 691
rect 672 552 696 691
rect 874 664 890 668
rect 911 663 930 668
rect 955 663 971 668
rect 278 546 304 550
rect 278 529 282 546
rect 299 529 304 546
rect 278 510 304 529
rect 278 493 282 510
rect 299 493 304 510
rect 278 484 304 493
rect 670 545 697 552
rect 670 528 676 545
rect 693 528 697 545
rect 670 509 697 528
rect 670 492 676 509
rect 693 492 697 509
rect 670 486 697 492
rect 279 400 303 484
rect 279 383 283 400
rect 300 383 303 400
rect 279 364 303 383
rect 279 347 283 364
rect 300 347 303 364
rect 279 223 303 347
rect 672 386 696 486
rect 672 369 676 386
rect 693 369 696 386
rect 917 377 930 379
rect 909 375 933 377
rect 672 350 696 369
rect 889 374 933 375
rect 889 357 912 374
rect 930 357 933 374
rect 889 356 933 357
rect 909 354 933 356
rect 919 350 930 354
rect 672 333 676 350
rect 693 333 696 350
rect 672 227 696 333
rect 671 224 697 227
rect 278 220 304 223
rect 671 195 697 198
rect 278 191 304 194
rect 279 41 303 191
rect 440 41 478 101
rect 672 41 696 195
<< via1 >>
rect 278 194 304 220
rect 671 198 697 224
<< metal2 >>
rect 0 617 763 635
rect 0 573 763 591
rect 0 463 763 481
rect 0 420 763 438
rect 0 293 762 311
rect 0 250 763 268
rect 668 224 700 225
rect 275 194 278 220
rect 304 219 307 220
rect 668 219 671 224
rect 304 201 671 219
rect 304 194 307 201
rect 668 198 671 201
rect 697 198 700 224
rect 668 196 700 198
rect 0 140 762 158
rect 0 98 760 115
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1634057701
transform 1 0 1040 0 -1 408
box 0 0 256 191
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1634057701
transform 1 0 1040 0 1 0
box 0 0 256 191
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1634057701
transform 1 0 1040 0 -1 732
box 0 0 256 191
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1634057701
transform 1 0 1040 0 1 323
box 0 0 256 191
use sky130_hilas_wellContact  sky130_hilas_wellContact_1
timestamp 1634057703
transform 1 0 1448 0 1 738
box 0 0 173 186
use sky130_hilas_wellContact  sky130_hilas_wellContact_0
timestamp 1634057703
transform 1 0 1851 0 1 731
box 0 0 173 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_0
timestamp 1634057705
transform 1 0 1332 0 1 436
box 0 0 223 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_2
timestamp 1634057705
transform 1 0 1332 0 1 760
box 0 0 223 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_1
timestamp 1634057705
transform 1 0 1332 0 1 575
box 0 0 223 186
use sky130_hilas_FGVaractorCapacitor  sky130_hilas_FGVaractorCapacitor_3
timestamp 1634057705
transform 1 0 1332 0 1 900
box 0 0 223 186
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_1
timestamp 1634057702
transform 1 0 1451 0 1 441
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_2
timestamp 1634057702
transform 1 0 1451 0 1 769
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_0
timestamp 1634057702
transform 1 0 1451 0 1 580
box 0 0 173 190
use sky130_hilas_TunCap01  sky130_hilas_TunCap01_3
timestamp 1634057702
transform 1 0 1451 0 1 900
box 0 0 173 190
<< labels >>
rlabel metal1 35 656 75 668 0 VTUN
port 1 nsew
rlabel metal1 955 663 971 668 0 VINJ
port 2 nsew
rlabel metal1 911 663 930 668 0 COLSEL1
port 3 nsew
rlabel metal1 874 664 890 668 0 COL1
port 4 nsew
rlabel metal1 440 658 478 668 0 GATE1
port 5 nsew
rlabel poly 642 279 659 294 0 FG3
rlabel metal1 279 663 303 668 0 VGND
port 14 nsew
rlabel metal1 672 663 696 668 0 VGND
port 14 nsew
rlabel metal1 672 63 696 69 0 VGND
port 14 nsew
rlabel metal1 279 63 303 69 0 VGND
port 14 nsew
rlabel metal1 440 63 478 72 0 GATE1
port 5 nsew
rlabel metal2 0 98 8 115 0 DRAIN4
port 15 nsew
rlabel metal2 0 140 6 158 0 ROW4
port 11 nsew
rlabel metal2 0 617 6 635 0 DRAIN1
port 16 nsew
rlabel metal2 0 573 6 591 0 ROW1
port 17 nsew
rlabel metal2 0 250 6 268 0 ROW3
port 18 nsew
rlabel metal2 0 293 6 311 0 DRAIN3
port 19 nsew
rlabel metal2 0 420 6 438 0 DRAIN2
port 20 nsew
rlabel metal2 0 463 6 481 0 ROW2
port 21 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
