magic
tech sky130A
timestamp 1627736296
<< psubdiff >>
rect -2715 816 2606 820
rect -2715 799 -2677 816
rect 2586 799 2606 816
rect -2715 796 2606 799
rect -2715 793 -2691 796
rect -2715 33 -2711 793
rect -2694 33 -2691 793
rect 2742 794 2766 820
rect -2715 17 -2691 33
rect 2742 85 2746 794
rect 2763 85 2766 794
rect 2742 65 2766 85
<< psubdiffcont >>
rect -2677 799 2586 816
rect -2711 33 -2694 793
rect 2746 85 2763 794
<< poly >>
rect -642 946 -593 968
rect -642 929 -632 946
rect -615 929 -593 946
rect -642 910 -593 929
rect -642 893 -632 910
rect -615 893 -593 910
rect -642 874 -593 893
rect -642 857 -632 874
rect -615 857 -593 874
rect 5 963 70 968
rect 5 946 43 963
rect 60 946 70 963
rect 5 929 70 946
rect 5 912 43 929
rect 60 912 70 929
rect 5 895 70 912
rect 5 878 43 895
rect 60 878 70 895
rect -642 833 -593 857
rect 5 861 70 878
rect 5 844 43 861
rect 60 844 70 861
rect 5 833 70 844
rect 2621 812 2727 818
rect 2621 795 2630 812
rect 2718 795 2727 812
rect 2621 790 2727 795
rect 2581 788 2727 790
rect -2682 772 2727 788
rect -2682 746 -2666 772
rect 2621 771 2727 772
rect -2682 730 2730 746
rect -2682 704 -2666 705
rect 2714 704 2730 730
rect -2682 688 2730 704
rect -2682 665 -2666 688
rect -2682 649 2730 665
rect 2714 624 2730 649
rect -2682 608 2730 624
rect -2682 586 -2666 608
rect -2682 570 2730 586
rect -2682 547 -2666 548
rect 2714 547 2730 570
rect -2682 531 2730 547
rect -2682 507 -2666 531
rect -2682 491 2730 507
rect -2682 469 -2666 470
rect 2714 469 2730 491
rect -2682 453 2730 469
rect -2682 427 -2666 453
rect -2682 411 2730 427
rect 2714 386 2730 411
rect -2682 370 2730 386
rect -2682 349 -2667 370
rect -2682 333 2730 349
rect 2714 311 2730 333
rect -2682 295 2730 311
rect -2682 273 -2666 295
rect -2682 257 2730 273
rect 2714 234 2730 257
rect -2682 218 2730 234
rect -2682 196 -2666 218
rect -2682 180 2730 196
rect 2714 158 2730 180
rect -2680 142 2730 158
rect -2680 121 -2664 142
rect -2680 105 2731 121
rect 2715 84 2731 105
rect -2677 68 2731 84
rect -2677 46 -2661 68
rect -2677 30 2730 46
rect 2714 7 2730 30
rect -62 -1 2730 7
rect -67 -18 -50 -1
rect -33 -18 -16 -1
rect 1 -18 18 -1
rect 35 -18 52 -1
rect 69 -18 86 -1
rect 103 -18 120 -1
rect 137 -9 2730 -1
rect 137 -18 174 -9
rect -62 -27 174 -18
<< polycont >>
rect -632 929 -615 946
rect -632 893 -615 910
rect -632 857 -615 874
rect 43 946 60 963
rect 43 912 60 929
rect 43 878 60 895
rect 43 844 60 861
rect 2630 795 2718 812
rect -50 -18 -33 -1
rect -16 -18 1 -1
rect 18 -18 35 -1
rect 52 -18 69 -1
rect 86 -18 103 -1
rect 120 -18 137 -1
<< npolyres >>
rect -593 868 5 968
<< locali >>
rect -635 964 -613 967
rect -635 947 -632 964
rect -615 947 -613 964
rect -635 946 -613 947
rect -635 929 -632 946
rect -615 929 -613 946
rect -635 928 -613 929
rect -635 911 -632 928
rect -615 911 -613 928
rect -635 910 -613 911
rect -635 893 -632 910
rect -615 893 -613 910
rect -635 892 -613 893
rect -635 875 -632 892
rect -615 875 -613 892
rect -635 874 -613 875
rect -635 857 -632 874
rect -615 857 -613 874
rect -635 856 -613 857
rect -635 855 -632 856
rect -640 839 -632 855
rect -615 855 -613 856
rect 39 963 63 971
rect 39 930 43 963
rect 60 930 63 963
rect 39 929 63 930
rect 39 912 43 929
rect 60 912 63 929
rect 39 911 63 912
rect 39 878 43 911
rect 60 878 63 911
rect 39 875 63 878
rect -615 839 -607 855
rect -640 836 -607 839
rect 39 844 43 875
rect 60 844 63 875
rect 39 836 63 844
rect -2711 799 -2677 816
rect 2586 812 2763 816
rect 2586 799 2630 812
rect -2711 795 2630 799
rect -2711 793 -2677 795
rect -2694 778 -2677 793
rect -287 789 601 795
rect -287 778 -277 789
rect -2694 776 -277 778
rect 592 778 601 789
rect 2718 794 2763 812
rect 2718 778 2746 794
rect 592 776 2746 778
rect 2746 68 2763 85
rect -2711 16 -2694 33
rect -33 -18 -30 -1
rect 1 -18 7 -1
rect 35 -18 43 -1
rect 69 -18 79 -1
rect 103 -18 115 -1
rect 137 -18 152 -1
<< viali >>
rect -632 947 -615 964
rect -632 911 -615 928
rect -632 875 -615 892
rect -632 839 -615 856
rect 43 946 60 947
rect 43 930 60 946
rect 43 895 60 911
rect 43 894 60 895
rect 43 861 60 875
rect 43 858 60 861
rect -2677 778 -287 795
rect 601 778 2718 795
rect -67 -18 -50 -1
rect -30 -18 -16 -1
rect -16 -18 -13 -1
rect 7 -18 18 -1
rect 18 -18 24 -1
rect 43 -18 52 -1
rect 52 -18 60 -1
rect 79 -18 86 -1
rect 86 -18 96 -1
rect 115 -18 120 -1
rect 120 -18 133 -1
rect 152 -18 169 -1
<< metal1 >>
rect -643 968 -402 1032
rect -641 964 -600 968
rect -641 947 -632 964
rect -615 947 -600 964
rect -641 928 -600 947
rect -641 911 -632 928
rect -615 911 -600 928
rect -641 892 -600 911
rect 32 947 73 979
rect 32 930 43 947
rect 60 930 73 947
rect 32 911 73 930
rect 32 902 43 911
rect -641 875 -632 892
rect -615 875 -600 892
rect -641 856 -600 875
rect -641 839 -632 856
rect -615 839 -600 856
rect -641 833 -600 839
rect 5 894 43 902
rect 60 894 73 911
rect 5 875 73 894
rect 5 858 43 875
rect 60 858 174 875
rect 5 832 174 858
rect -2716 814 -279 816
rect -2722 810 -279 814
rect -2722 795 -2667 810
rect -2722 778 -2677 795
rect -287 778 -279 810
rect -2722 775 -279 778
rect -2722 -50 -2681 775
rect -62 25 174 832
rect 601 815 2737 816
rect 595 810 2737 815
rect 595 778 601 810
rect 2687 795 2737 810
rect 2718 778 2737 795
rect 595 776 2737 778
rect 595 775 2721 776
rect -74 -1 174 25
rect -74 -18 -67 -1
rect -50 -18 -30 -1
rect -13 -18 7 -1
rect 24 -18 43 -1
rect 60 -18 79 -1
rect 96 -18 115 -1
rect 133 -18 152 -1
rect 169 -18 174 -1
rect -74 -57 174 -18
<< via1 >>
rect -2667 795 -287 810
rect -2667 784 -287 795
rect 601 795 2687 810
rect 601 784 2687 795
<< metal2 >>
rect -2749 810 2798 820
rect -2749 784 -2667 810
rect -287 784 601 810
rect 2687 784 2798 810
rect -2749 681 2798 784
rect -2749 51 2798 191
<< labels >>
rlabel metal1 -642 983 -404 1022 0 INPUT
port 2 nsew
rlabel metal1 -74 -57 174 -30 0 OUTPUT
port 3 nsew
rlabel metal1 -2722 -50 -2681 -39 0 VGND
port 4 nsew
<< end >>
