* Copyright 2020 The Hilas PDK Authors
* 
* This file is part of HILAS.
* 
* HILAS is free software: you can redistribute it and/or modify
* it under the terms of the GNU Lesser General Public License as published by
* the Free Software Foundation, version 3 of the License.
* 
* HILAS is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU Lesser General Public License for more details.
* 
* You should have received a copy of the GNU Lesser General Public License
* along with HILAS.  If not, see <https://www.gnu.org/licenses/>.
* 
* Licensed under the Lesser General Public License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
* https://www.gnu.org/licenses/lgpl-3.0.en.html
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* 
* SPDX-License-Identifier: LGPL-3.0
* 
* 

* NGSPICE file created from sky130_hilas_Tgate4Double01.ext - technology: sky130A

.subckt sky130_hilas_TgateDouble01 a_n40_n314# $SUB a_n468_n112# output w_n502_n362#
+ a_290_n314#
X0 a_n196_n192# a_n468_n112# w_n502_n362# w_n502_n362# sky130_fd_pr__pfet_01v8 w=320000u l=400000u
X1 $SUB a_n468_n112# a_n196_n192# $SUB sky130_fd_pr__nfet_01v8 w=300000u l=400000u
X2 output a_n468_n112# a_n40_n314# $SUB sky130_fd_pr__nfet_01v8 w=310000u l=400000u
X3 output a_n468_n112# a_290_n314# w_n502_n362# sky130_fd_pr__pfet_01v8 w=310000u l=400000u
X4 output a_n196_n192# a_n40_n314# w_n502_n362# sky130_fd_pr__pfet_01v8 w=310000u l=400000u
X5 output a_n196_n192# a_290_n314# $SUB sky130_fd_pr__nfet_01v8 w=310000u l=400000u
.ends

.subckt sky130_hilas_Tgate4Double01 VPWR INPUT1_1 INPUT2_1 SELECT1 SELECT2 INPUT2_2
+ INPUT1_2 SELECT3 INPUT2_3 SELECT4 INPUT2_4 INPUT1_4 OUTPUT4 OUTPUT3 OUTPUT2 OUTPUT1
Xsky130_hilas_TgateDouble01_0 INPUT1_1 VPWR SELECT1 OUTPUT1 VPWR INPUT2_1 sky130_hilas_TgateDouble01
Xsky130_hilas_TgateDouble01_1 INPUT1_4 VPWR SELECT4 OUTPUT4 VPWR INPUT2_4 sky130_hilas_TgateDouble01
Xsky130_hilas_TgateDouble01_2 Input1_3 VPWR SELECT3 OUTPUT3 VPWR INPUT2_3 sky130_hilas_TgateDouble01
Xsky130_hilas_TgateDouble01_3 INPUT1_2 VPWR SELECT2 OUTPUT2 VPWR INPUT2_2 sky130_hilas_TgateDouble01
.ends

