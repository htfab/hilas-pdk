VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_pFETLarge
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pFETLarge ;
  ORIGIN -0.640 -4.190 ;
  SIZE 4.640 BY 5.990 ;
  PIN Gate
    PORT
      LAYER met2 ;
        RECT 0.640 4.200 0.960 5.020 ;
    END
  END Gate
  PIN Source
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 0.880 5.320 1.200 9.790 ;
    END
  END Source
  PIN Drain
    USE ANALOG ;
    PORT
      LAYER met2 ;
        RECT 4.660 4.650 5.010 9.080 ;
    END
  END Drain
  PIN Well
    USE ANALOG ;
    PORT
      LAYER met1 ;
        RECT 4.780 9.870 5.040 10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.780 4.190 5.040 9.360 ;
    END
  END Well
  OBS
      LAYER li1 ;
        RECT 0.830 4.200 5.060 9.870 ;
      LAYER met1 ;
        RECT 0.930 4.200 4.500 9.980 ;
      LAYER met2 ;
        RECT 1.480 9.360 4.780 9.800 ;
        RECT 1.480 5.040 4.380 9.360 ;
        RECT 1.240 4.370 4.380 5.040 ;
        RECT 1.240 4.200 4.780 4.370 ;
  END
END sky130_hilas_pFETLarge
END LIBRARY

