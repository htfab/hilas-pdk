magic
tech sky130A
timestamp 1634057768
<< metal3 >>
rect 0 0 230 228
<< mimcap >>
rect 15 111 215 214
rect 15 98 100 111
rect 114 98 215 111
rect 15 14 215 98
<< mimcapcontact >>
rect 100 98 114 111
<< metal4 >>
rect 85 123 130 124
rect 83 111 135 123
rect 83 98 100 111
rect 114 98 135 111
rect 83 74 135 98
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
