magic
tech sky130A
timestamp 1628616752
<< checkpaint >>
rect 2429 2713 6381 2754
rect 2429 2700 6489 2713
rect 322 2251 6489 2700
rect -1299 2115 6489 2251
rect -1299 -58 6491 2115
rect -1296 -591 6491 -58
rect -1296 -630 6157 -591
rect -1296 -652 3987 -630
rect -1296 -656 3210 -652
<< error_s >>
rect 413 1136 419 1142
rect 518 1136 524 1142
rect 1384 1136 1390 1142
rect 1489 1136 1495 1142
rect 2463 1136 2469 1142
rect 2568 1136 2574 1142
rect 839 1126 845 1132
rect 892 1126 898 1132
rect 1010 1126 1016 1132
rect 1063 1126 1069 1132
rect 2889 1126 2895 1132
rect 2942 1126 2948 1132
rect 407 1072 413 1078
rect 524 1072 530 1078
rect 833 1076 839 1082
rect 898 1076 904 1082
rect 1004 1076 1010 1082
rect 1069 1076 1075 1082
rect 1378 1072 1384 1078
rect 1495 1072 1501 1078
rect 2457 1072 2463 1078
rect 2574 1072 2580 1078
rect 2883 1076 2889 1082
rect 2948 1076 2954 1082
rect 413 1019 419 1025
rect 518 1019 524 1025
rect 839 1017 845 1023
rect 892 1017 898 1023
rect 1010 1017 1016 1023
rect 1063 1017 1069 1023
rect 1384 1019 1390 1025
rect 1489 1019 1495 1025
rect 2463 1019 2469 1025
rect 2568 1019 2574 1025
rect 2889 1017 2895 1023
rect 2942 1017 2948 1023
rect 833 967 839 973
rect 898 967 904 973
rect 1004 967 1010 973
rect 1069 967 1075 973
rect 2883 967 2889 973
rect 2948 967 2954 973
rect 182 959 195 964
rect 196 959 209 963
rect 182 956 209 959
rect 407 955 413 961
rect 524 955 530 961
rect 1378 955 1384 961
rect 1495 955 1501 961
rect 1699 959 1712 963
rect 1713 959 1726 964
rect 1699 956 1726 959
rect 2457 955 2463 961
rect 2574 955 2580 961
rect 413 834 419 840
rect 518 834 524 840
rect 1384 834 1390 840
rect 1489 834 1495 840
rect 2463 834 2469 840
rect 2568 834 2574 840
rect 839 828 845 834
rect 892 828 898 834
rect 1010 828 1016 834
rect 1063 828 1069 834
rect 2889 828 2895 834
rect 2942 828 2948 834
rect 833 778 839 784
rect 898 778 904 784
rect 1004 778 1010 784
rect 1069 778 1075 784
rect 2883 778 2889 784
rect 2948 778 2954 784
rect 407 770 413 776
rect 524 770 530 776
rect 1378 770 1384 776
rect 1495 770 1501 776
rect 2457 770 2463 776
rect 2574 770 2580 776
rect 413 718 419 724
rect 518 718 524 724
rect 1384 718 1390 724
rect 1489 718 1495 724
rect 839 711 845 717
rect 892 711 898 717
rect 1010 711 1016 717
rect 1063 711 1069 717
rect 1924 715 1925 727
rect 2463 718 2469 724
rect 2568 718 2574 724
rect 1938 701 1939 713
rect 2889 711 2895 717
rect 2942 711 2948 717
rect 833 661 839 667
rect 898 661 904 667
rect 1004 661 1010 667
rect 1069 661 1075 667
rect 2883 661 2889 667
rect 2948 661 2954 667
rect 407 654 413 660
rect 524 654 530 660
rect 1378 654 1384 660
rect 1495 654 1501 660
rect 2457 654 2463 660
rect 2574 654 2580 660
rect 87 614 89 622
rect 2137 614 2138 622
rect 0 601 1 609
rect 81 601 82 609
rect 1843 603 1844 609
rect 1843 595 1845 603
rect 1924 601 1925 609
rect 416 538 422 544
rect 521 538 527 544
rect 1387 538 1393 544
rect 1492 538 1498 544
rect 2465 538 2471 544
rect 2570 538 2576 544
rect 842 528 848 534
rect 895 528 901 534
rect 1013 528 1019 534
rect 1066 528 1072 534
rect 2891 528 2897 534
rect 2944 528 2950 534
rect 410 474 416 480
rect 527 474 533 480
rect 836 478 842 484
rect 901 478 907 484
rect 1007 478 1013 484
rect 1072 478 1078 484
rect 1381 474 1387 480
rect 1498 474 1504 480
rect 2459 474 2465 480
rect 2576 474 2582 480
rect 2885 478 2891 484
rect 2950 478 2956 484
rect 416 421 422 427
rect 521 421 527 427
rect 842 419 848 425
rect 895 419 901 425
rect 1013 419 1019 425
rect 1066 419 1072 425
rect 1387 421 1393 427
rect 1492 421 1498 427
rect 2465 421 2471 427
rect 2570 421 2576 427
rect 2891 419 2897 425
rect 2944 419 2950 425
rect 836 369 842 375
rect 901 369 907 375
rect 1007 369 1013 375
rect 1072 369 1078 375
rect 2885 369 2891 375
rect 2950 369 2956 375
rect 185 361 198 366
rect 199 361 212 365
rect 185 358 212 361
rect 410 357 416 363
rect 527 357 533 363
rect 1381 357 1387 363
rect 1498 357 1504 363
rect 1702 361 1715 365
rect 1716 361 1729 366
rect 1702 358 1729 361
rect 2459 357 2465 363
rect 2576 357 2582 363
rect 416 236 422 242
rect 521 236 527 242
rect 1387 236 1393 242
rect 1492 236 1498 242
rect 2465 236 2471 242
rect 2570 236 2576 242
rect 842 230 848 236
rect 895 230 901 236
rect 1013 230 1019 236
rect 1066 230 1072 236
rect 2891 230 2897 236
rect 2944 230 2950 236
rect 836 180 842 186
rect 901 180 907 186
rect 1007 180 1013 186
rect 1072 180 1078 186
rect 2885 180 2891 186
rect 2950 180 2956 186
rect 410 172 416 178
rect 527 172 533 178
rect 1381 172 1387 178
rect 1498 172 1504 178
rect 2459 172 2465 178
rect 2576 172 2582 178
rect 416 120 422 126
rect 521 120 527 126
rect 1387 120 1393 126
rect 1492 120 1498 126
rect 842 113 848 119
rect 895 113 901 119
rect 1013 113 1019 119
rect 1066 113 1072 119
rect 1926 117 1928 129
rect 2465 120 2471 126
rect 2570 120 2576 126
rect 1926 69 1927 117
rect 1940 103 1942 115
rect 2891 113 2897 119
rect 2944 113 2950 119
rect 1940 83 1941 103
rect 836 63 842 69
rect 901 63 907 69
rect 1007 63 1013 69
rect 1072 63 1078 69
rect 2885 63 2891 69
rect 2950 63 2956 69
rect 410 56 416 62
rect 527 56 533 62
rect 1381 56 1387 62
rect 1498 56 1504 62
rect 2459 56 2465 62
rect 2576 56 2582 62
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_1
timestamp 1628616734
transform 1 0 3059 0 1 637
box 0 0 2692 1487
use sky130_hilas_WTA4Stage01  sky130_hilas_WTA4Stage01_0
timestamp 1628616734
transform 1 0 3061 0 1 39
box 0 0 2692 1487
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_1
timestamp 1628616737
transform 1 0 952 0 1 598
box 0 0 4572 1472
use sky130_hilas_swc4x2cell  sky130_hilas_swc4x2cell_0
timestamp 1628616737
transform 1 0 955 0 1 0
box 0 0 4572 1472
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
