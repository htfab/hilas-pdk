magic
tech sky130A
timestamp 1628704408
<< error_s >>
rect 65 660 115 666
rect 388 661 438 667
rect 545 660 573 667
rect 687 661 715 667
rect 65 618 115 624
rect 388 619 438 625
rect 545 618 573 625
rect 687 619 715 625
rect 136 594 186 600
rect 316 589 367 595
rect 496 589 524 595
rect 736 589 764 595
rect 136 552 186 558
rect 316 547 367 553
rect 496 547 524 553
rect 736 547 764 553
rect 65 485 115 491
rect 388 486 438 492
rect 545 485 573 492
rect 687 486 715 492
rect 65 443 115 449
rect 388 444 438 450
rect 545 443 573 450
rect 687 444 715 450
rect 136 419 186 425
rect 316 414 367 420
rect 496 414 524 420
rect 736 414 764 420
rect 136 377 186 383
rect 316 372 367 378
rect 496 372 524 378
rect 736 372 764 378
rect 65 310 115 316
rect 388 311 438 317
rect 545 310 573 317
rect 687 311 715 317
rect 65 268 115 274
rect 388 269 438 275
rect 545 268 573 275
rect 687 269 715 275
rect 136 244 186 250
rect 316 239 367 245
rect 496 239 524 245
rect 736 239 764 245
rect 136 202 186 208
rect 316 197 367 203
rect 496 197 524 203
rect 736 197 764 203
rect 65 135 115 141
rect 388 136 438 142
rect 545 135 573 142
rect 687 136 715 142
rect 65 93 115 99
rect 388 94 438 100
rect 545 93 573 100
rect 687 94 715 100
rect 136 69 186 75
rect 316 64 367 70
rect 496 64 524 70
rect 736 64 764 70
rect 136 27 186 33
rect 316 22 367 28
rect 496 22 524 28
rect 736 22 764 28
<< nwell >>
rect 0 576 11 596
<< metal1 >>
rect 34 691 63 700
rect 465 694 496 700
rect 766 695 790 700
rect 34 0 63 12
rect 465 0 496 6
rect 766 0 790 5
<< metal2 >>
rect 0 636 16 656
rect 860 543 870 575
rect 0 461 17 481
rect 860 368 870 400
rect 0 286 19 306
rect 860 193 870 225
rect 0 111 16 131
rect 860 18 870 50
use sky130_hilas_StepUpDigital  StepUpDigital_2
timestamp 1628704371
transform 1 0 -19 0 1 569
box 0 0 870 175
use sky130_hilas_StepUpDigital  StepUpDigital_1
timestamp 1628704371
transform 1 0 -19 0 1 394
box 0 0 870 175
use sky130_hilas_StepUpDigital  StepUpDigital_3
timestamp 1628704371
transform 1 0 -19 0 1 44
box 0 0 870 175
use sky130_hilas_StepUpDigital  StepUpDigital_0
timestamp 1628704371
transform 1 0 -19 0 1 219
box 0 0 870 175
<< labels >>
rlabel metal1 34 4 63 9 0 VINJ
port 6 nsew
rlabel metal2 0 111 11 131 0 OUTPUT4
port 10 nsew
rlabel metal2 860 543 870 575 0 INPUT1
port 12 nsew
rlabel metal2 860 368 870 400 0 INPUT2
port 13 nsew
rlabel metal2 860 193 870 225 0 INPUT3
port 14 nsew
rlabel metal2 860 18 870 50 0 INPUT4
port 15 nsew
rlabel metal2 0 286 8 306 0 OUTPUT3
port 9 nsew
rlabel metal2 0 461 7 481 0 OUTPUT2
port 8 nsew
rlabel metal2 0 636 7 656 0 OUTPUT1
port 7 nsew
rlabel metal1 465 0 496 6 0 VGND
port 11 nsew
rlabel metal1 465 694 496 700 0 VGND
port 11 nsew
rlabel metal1 34 691 63 700 0 VINJ
port 6 nsew
rlabel metal1 766 695 790 700 0 VPWR
port 5 nsew
rlabel metal1 766 0 790 5 0 VPWR
port 5 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
