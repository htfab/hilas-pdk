magic
tech sky130A
magscale 1 2
timestamp 1632255311
<< error_s >>
rect 302 1592 380 1598
rect 624 1592 702 1598
rect 946 1592 1024 1598
rect 302 1508 380 1514
rect 624 1508 702 1514
rect 946 1508 1024 1514
rect 1222 1446 1466 1638
rect 1478 1446 1720 1638
rect 1912 1592 1990 1598
rect 2234 1592 2312 1598
rect 2556 1592 2634 1598
rect 2878 1592 2956 1598
rect 3200 1592 3278 1598
rect 1810 1468 1822 1540
rect 1912 1508 1990 1514
rect 2234 1508 2312 1514
rect 2556 1508 2634 1514
rect 2878 1508 2956 1514
rect 3200 1508 3278 1514
rect 1476 1426 1720 1446
rect 302 1400 380 1406
rect 620 1400 698 1406
rect 942 1400 1020 1406
rect 1264 1400 1342 1406
rect 1434 1396 1720 1426
rect 1908 1400 1986 1406
rect 2230 1400 2308 1406
rect 2552 1400 2630 1406
rect 2874 1400 2952 1406
rect 3200 1400 3278 1406
rect 1476 1362 1718 1396
rect 302 1316 380 1322
rect 362 1276 450 1280
rect 520 1276 522 1348
rect 1476 1322 1730 1362
rect 620 1316 698 1322
rect 942 1316 1020 1322
rect 1264 1316 1342 1322
rect 1476 1316 1738 1322
rect 1002 1276 1090 1280
rect 302 1208 380 1214
rect 404 1208 422 1238
rect 620 1208 698 1214
rect 942 1208 1020 1214
rect 1044 1208 1062 1238
rect 389 1193 432 1208
rect 1029 1193 1074 1208
rect 404 1172 432 1193
rect 1044 1172 1074 1193
rect 354 1130 380 1162
rect 417 1157 432 1172
rect 381 1130 432 1135
rect 302 1124 380 1130
rect 354 1120 380 1124
rect 396 1114 422 1120
rect 520 1084 522 1156
rect 620 1124 698 1130
rect 722 1044 740 1082
rect 750 1063 768 1094
rect 842 1084 848 1138
rect 998 1130 1020 1162
rect 1059 1157 1074 1172
rect 1222 1158 1464 1316
rect 1476 1204 1786 1316
rect 1808 1276 1818 1348
rect 1908 1316 1986 1322
rect 2230 1316 2308 1322
rect 2552 1316 2630 1322
rect 2874 1316 2952 1322
rect 1970 1276 2056 1282
rect 2292 1276 2378 1282
rect 1908 1208 1986 1214
rect 2012 1208 2028 1240
rect 2230 1208 2308 1214
rect 2334 1208 2350 1240
rect 3034 1234 3052 1276
rect 2552 1208 2630 1214
rect 2874 1208 2952 1214
rect 1488 1184 1786 1204
rect 1808 1192 1832 1204
rect 1997 1193 2040 1208
rect 2319 1196 2362 1208
rect 2319 1193 2394 1196
rect 1488 1172 1790 1184
rect 1488 1158 1786 1172
rect 1025 1130 1074 1135
rect 942 1124 1020 1130
rect 998 1120 1020 1124
rect 1222 1120 1786 1158
rect 1790 1150 1792 1158
rect 1808 1128 1834 1192
rect 2012 1174 2040 1193
rect 2334 1190 2394 1193
rect 2334 1184 2400 1190
rect 2334 1174 2362 1184
rect 1964 1130 1986 1166
rect 2025 1159 2040 1174
rect 2347 1168 2362 1174
rect 1991 1130 2040 1139
rect 2286 1130 2308 1164
rect 2342 1156 2372 1168
rect 2724 1140 2730 1170
rect 2794 1142 2796 1180
rect 2313 1130 2362 1137
rect 2828 1136 2830 1202
rect 1790 1120 1792 1128
rect 1040 1114 1062 1120
rect 1222 1112 1792 1120
rect 750 1046 790 1063
rect 1222 1062 1644 1112
rect 1762 1100 1792 1112
rect 1808 1120 1832 1128
rect 1908 1124 1986 1130
rect 2230 1124 2308 1130
rect 2552 1124 2630 1130
rect 2874 1124 2952 1130
rect 1808 1114 1838 1120
rect 2006 1114 2028 1124
rect 2286 1122 2308 1124
rect 2328 1114 2350 1122
rect 1808 1108 1900 1114
rect 1808 1084 2028 1108
rect 750 1044 768 1046
rect 720 1042 778 1044
rect 1434 1042 1442 1062
rect 302 1016 380 1022
rect 620 1016 698 1022
rect 722 1016 740 1042
rect 750 1030 768 1042
rect 942 1016 1020 1022
rect 1264 1016 1342 1022
rect 722 1015 752 1016
rect 722 1010 740 1015
rect 710 1008 744 1010
rect 722 1002 740 1008
rect 1464 1004 1718 1062
rect 1908 1040 1986 1046
rect 1804 1012 1846 1038
rect 1854 1028 1889 1040
rect 1854 1025 1873 1028
rect 1854 1012 1858 1025
rect 2608 1022 2632 1044
rect 3034 1042 3052 1084
rect 2230 1016 2308 1022
rect 2552 1016 2632 1022
rect 2874 1016 2952 1022
rect 1854 1004 1869 1012
rect 2608 1004 2632 1016
rect 2642 1004 2666 1010
rect 302 932 380 938
rect 520 892 522 964
rect 620 932 698 938
rect 942 932 1020 938
rect 1264 932 1342 938
rect 1434 860 1442 892
rect 1476 860 1718 990
rect 1770 978 1880 1004
rect 1908 956 1986 962
rect 2116 958 2184 960
rect 2054 926 2086 946
rect 2176 938 2193 957
rect 2828 944 2862 966
rect 2230 932 2308 938
rect 2552 932 2630 938
rect 2874 932 2952 938
rect 2096 924 2150 926
rect 2096 874 2128 924
rect 2862 910 2896 932
rect 3034 860 3052 892
rect 3076 860 3328 1396
rect 178 628 1464 860
rect 1476 628 3074 860
rect 3076 628 3398 860
rect 302 560 380 566
rect 624 560 702 566
rect 946 560 1024 566
rect 1268 560 1346 566
rect 302 476 380 482
rect 624 476 702 482
rect 946 476 1024 482
rect 1268 476 1346 482
rect 1478 436 1720 606
rect 1912 560 1990 566
rect 2234 560 2312 566
rect 2556 560 2634 566
rect 2878 560 2956 566
rect 3200 560 3278 566
rect 1810 436 1822 508
rect 1912 476 1990 482
rect 2234 476 2312 482
rect 2556 476 2634 482
rect 2878 476 2956 482
rect 3200 476 3278 482
<< nwell >>
rect 474 990 2760 1004
<< poly >>
rect 396 1114 448 1120
rect 1040 1114 1092 1120
rect 1362 1114 1414 1122
rect 1684 1114 1736 1120
rect 2006 1114 2058 1124
rect 2328 1114 2380 1122
<< locali >>
rect 796 1004 830 1006
rect 2590 1004 2632 1160
rect 2724 1004 2758 1140
rect 474 958 2760 1004
rect 474 246 508 958
rect 606 0 640 892
rect 796 246 830 958
rect 932 0 966 884
rect 1114 246 1148 958
rect 1252 0 1286 900
rect 1438 246 1472 958
rect 1576 0 1610 890
rect 1762 250 1796 958
rect 1896 0 1930 900
rect 2082 252 2116 958
rect 2220 0 2254 900
rect 2404 250 2438 958
rect 2540 0 2574 896
rect 2726 244 2760 958
rect 2862 0 2896 932
<< metal1 >>
rect 1348 710 2038 744
rect 1658 204 1694 512
rect 1998 342 2038 710
rect 608 0 3316 46
<< metal2 >>
rect 0 1154 1410 1192
rect 0 1150 58 1154
rect 0 990 412 1002
rect 696 990 740 1082
rect 1680 992 1730 1144
rect 1680 990 1736 992
rect 0 960 1736 990
rect 52 912 92 960
rect 380 930 1736 960
rect 2022 616 2062 1136
rect 0 574 2062 616
rect 2342 420 2372 1168
rect 2542 1136 2774 1192
rect 2692 1134 2774 1136
rect 0 380 2374 420
rect 0 378 28 380
rect 0 156 1708 196
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_9
timestamp 1632251409
transform 1 0 62 0 1 1128
box 0 0 66 110
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_11
timestamp 1632251409
transform 1 0 62 0 1 676
box 0 0 66 110
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_12
timestamp 1632251409
transform 1 0 62 0 1 488
box 0 0 66 110
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_10
timestamp 1632251409
transform 1 0 58 0 1 866
box 0 0 66 110
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_8
timestamp 1632251409
transform 1 0 404 0 1 1136
box 0 0 66 110
use sky130_hilas_DAC6TransistorStack01a  sky130_hilas_DAC6TransistorStack01a_0
timestamp 1632255311
transform 1 0 18 0 1 352
box 160 84 504 1286
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_7
timestamp 1632251409
transform 0 1 704 -1 0 1096
box 0 0 66 110
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_6
timestamp 1632251409
transform 1 0 1044 0 1 1136
box 0 0 66 110
use sky130_hilas_li2m1  sky130_hilas_li2m1_6
timestamp 1632251332
transform 1 0 946 0 1 14
box 0 0 46 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_0
timestamp 1632251332
transform 1 0 622 0 1 14
box 0 0 46 58
use sky130_hilas_DAC6TransistorStack01  sky130_hilas_DAC6TransistorStack01_0
array 0 2 322 0 0 1132
timestamp 1632255311
transform 1 0 340 0 1 352
box 158 84 504 1286
use sky130_hilas_DAC6TransistorStack01b  sky130_hilas_DAC6TransistorStack01b_0
timestamp 1632255311
transform 1 0 1306 0 1 352
box 170 84 552 1286
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_5
timestamp 1632251409
transform 1 0 1366 0 1 1138
box 0 0 66 110
use sky130_hilas_li2m1  sky130_hilas_li2m1_7
timestamp 1632251332
transform 1 0 1266 0 1 14
box 0 0 46 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_1
timestamp 1632251332
transform 1 0 1590 0 1 14
box 0 0 46 58
use sky130_hilas_DAC6TransistorStack01c  sky130_hilas_DAC6TransistorStack01c_0
timestamp 1632255311
transform 1 0 1628 0 1 352
box 158 84 534 1286
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_3
timestamp 1632251409
transform 1 0 2012 0 1 1138
box 0 0 66 110
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_4
timestamp 1632251409
transform 1 0 1690 0 1 1136
box 0 0 66 110
use sky130_hilas_li2m1  sky130_hilas_li2m1_5
timestamp 1632251332
transform 1 0 1910 0 1 14
box 0 0 46 58
use sky130_hilas_m12m2  sky130_hilas_m12m2_0
timestamp 1632251372
transform 1 0 1670 0 1 164
box 0 0 64 64
use sky130_hilas_DAC6TransistorStack01  sky130_hilas_DAC6TransistorStack01_2
array 0 2 322 0 0 1132
timestamp 1632255311
transform 1 0 1950 0 1 352
box 158 84 504 1286
use sky130_hilas_poly2m2  sky130_hilas_poly2m2_2
timestamp 1632251409
transform 1 0 2334 0 1 1138
box 0 0 66 110
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632251356
transform 1 0 2728 0 1 1130
box 0 0 68 66
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1632251356
transform 1 0 2594 0 1 1130
box 0 0 68 66
use sky130_hilas_li2m1  sky130_hilas_li2m1_2
timestamp 1632251332
transform 1 0 2234 0 1 14
box 0 0 46 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_4
timestamp 1632251332
transform 1 0 2876 0 1 14
box 0 0 46 58
use sky130_hilas_li2m1  sky130_hilas_li2m1_3
timestamp 1632251332
transform 1 0 2554 0 1 14
box 0 0 46 58
use sky130_hilas_DAC6TransistorStack01a  sky130_hilas_DAC6TransistorStack01a_1
timestamp 1632255311
transform 1 0 2916 0 1 352
box 160 84 504 1286
<< labels >>
rlabel metal2 2 1150 22 1192 0 A4
port 5 nsew analog default
rlabel metal2 0 960 20 1002 0 A3
port 4 nsew analog default
rlabel metal2 2 574 22 616 0 A2
port 3 nsew analog default
rlabel metal2 2 378 22 420 0 A1
port 2 nsew analog default
rlabel metal2 0 156 16 196 0 A0
port 1 nsew analog default
rlabel metal2 2542 1164 2692 1192 0 VPWR
port 6 nsew analog default
rlabel metal1 3292 0 3316 46 0 OUT
port 7 nsew analog default
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
