magic
tech sky130A
timestamp 1632494644
<< nwell >>
rect -289 41 -33 232
<< mvpmos >>
rect -222 126 -172 180
<< mvpdiff >>
rect -251 174 -222 180
rect -251 132 -247 174
rect -229 132 -222 174
rect -251 126 -222 132
rect -172 169 -142 180
rect -172 152 -166 169
rect -147 152 -142 169
rect -172 126 -142 152
<< mvpdiffc >>
rect -247 132 -229 174
rect -166 152 -147 169
<< nsubdiff >>
rect -142 169 -97 180
rect -142 152 -128 169
rect -109 152 -97 169
rect -142 125 -97 152
<< nsubdiffcont >>
rect -128 152 -109 169
<< poly >>
rect -222 180 -172 193
rect -222 117 -172 126
rect -289 100 -172 117
<< locali >>
rect -255 174 -221 176
rect -255 132 -247 174
rect -229 132 -221 174
rect -166 169 -106 177
rect -147 152 -128 169
rect -109 152 -106 169
rect -166 138 -106 152
rect -166 121 -165 138
rect -148 121 -127 138
rect -110 121 -106 138
rect -166 117 -106 121
<< viali >>
rect -165 121 -148 138
rect -127 121 -110 138
<< metal1 >>
rect -166 194 -150 232
rect -166 141 -107 194
rect -168 138 -107 141
rect -168 121 -165 138
rect -148 121 -127 138
rect -110 121 -107 138
rect -168 117 -107 121
rect -166 115 -107 117
rect -166 42 -150 115
<< metal2 >>
rect -289 140 -280 158
rect -250 140 -33 158
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1632488964
transform 1 0 -266 0 -1 156
box -14 -15 20 18
<< end >>
