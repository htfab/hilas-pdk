magic
tech sky130A
timestamp 1634057852
<< checkpaint >>
rect -630 -517 1035 1121
<< psubdiff >>
rect 398 31 399 114
<< locali >>
rect 373 490 392 579
rect 373 25 399 114
<< metal1 >>
rect 68 541 103 604
rect 68 525 330 541
rect 364 550 471 604
rect 364 541 383 550
rect 356 525 383 541
rect 68 524 383 525
rect 409 524 471 550
rect 68 510 471 524
rect 68 509 383 510
rect 68 483 328 509
rect 354 484 383 509
rect 409 484 471 510
rect 354 483 471 484
rect 68 473 471 483
rect 68 419 471 442
rect 68 392 119 419
rect 146 392 174 419
rect 201 392 471 419
rect 68 362 471 392
rect 68 361 174 362
rect 68 334 118 361
rect 145 335 174 361
rect 201 335 471 362
rect 145 334 471 335
rect 68 278 471 334
rect 68 277 174 278
rect 68 250 119 277
rect 146 251 174 277
rect 201 251 471 278
rect 146 250 471 251
rect 68 227 471 250
rect 68 200 119 227
rect 146 225 471 227
rect 146 200 172 225
rect 68 198 172 200
rect 199 198 471 225
rect 68 163 471 198
rect 68 100 471 127
rect 68 74 344 100
rect 370 74 392 100
rect 418 74 471 100
rect 68 59 471 74
rect 68 33 342 59
rect 368 33 391 59
rect 417 33 471 59
rect 68 3 471 33
rect 68 0 104 3
rect 373 1 471 3
rect 372 0 471 1
<< via1 >>
rect 330 525 356 551
rect 383 524 409 550
rect 328 483 354 509
rect 383 484 409 510
rect 119 392 146 419
rect 174 392 201 419
rect 118 334 145 361
rect 174 335 201 362
rect 119 250 146 277
rect 174 251 201 278
rect 119 200 146 227
rect 172 198 199 225
rect 344 74 370 100
rect 392 74 418 100
rect 342 33 368 59
rect 391 33 417 59
<< metal2 >>
rect 104 419 234 604
rect 104 392 119 419
rect 146 392 174 419
rect 201 392 234 419
rect 104 362 234 392
rect 104 361 174 362
rect 104 334 118 361
rect 145 335 174 361
rect 201 335 234 362
rect 145 334 234 335
rect 104 278 234 334
rect 104 277 174 278
rect 104 250 119 277
rect 146 251 174 277
rect 201 251 234 278
rect 146 250 234 251
rect 104 227 234 250
rect 104 200 119 227
rect 146 225 234 227
rect 146 200 172 225
rect 104 198 172 200
rect 199 198 234 225
rect 104 0 234 198
rect 312 551 442 604
rect 312 525 330 551
rect 356 550 442 551
rect 356 525 383 550
rect 312 524 383 525
rect 409 524 442 550
rect 312 510 442 524
rect 312 509 383 510
rect 312 483 328 509
rect 354 484 383 509
rect 409 484 442 510
rect 354 483 442 484
rect 312 462 442 483
rect 312 132 441 462
rect 312 100 442 132
rect 312 74 344 100
rect 370 74 392 100
rect 418 74 442 100
rect 312 59 442 74
rect 312 33 342 59
rect 368 33 391 59
rect 417 33 442 59
rect 312 0 442 33
use sky130_hilas_DecoupVinj00  CapDeco_1
timestamp 1634057788
transform 1 0 0 0 1 113
box 0 0 405 307
use sky130_hilas_DecoupVinj00  CapDeco_0
timestamp 1634057788
transform 1 0 0 0 -1 491
box 0 0 405 307
<< labels >>
rlabel metal1 82 0 91 63 0 VGND 
port 1 nsew
rlabel metal1 456 0 471 63 0 VGND 
port 1 nsew
rlabel metal2 104 594 234 604 0 VINJ
port 1 nsew
rlabel metal2 312 596 442 604 0 VGND
port 2 nsew
rlabel metal2 104 0 234 12 0 VINJ
port 1 nsew
rlabel metal2 312 0 442 12 0 VGND
port 2 nsew
rlabel metal1 454 256 471 350 0 VINJ
port 1 nsew
rlabel metal1 68 254 85 350 0 VINJ
port 1 nsew
rlabel metal1 82 541 90 604 0 VGND
port 3 nsew
rlabel metal1 461 541 471 604 0 VGND
port 2 nsew
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
