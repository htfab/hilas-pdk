magic
tech sky130A
timestamp 1634057701
<< checkpaint >>
rect -607 -603 687 745
<< error_s >>
rect 67 139 117 145
rect 67 97 117 103
rect 67 70 117 76
rect 139 70 189 76
rect 67 28 117 34
rect 139 28 189 34
<< nwell >>
rect 0 0 256 191
<< mvpmos >>
rect 67 103 117 139
rect 67 34 117 70
rect 139 34 189 70
<< mvpdiff >>
rect 38 126 67 139
rect 38 109 42 126
rect 60 109 67 126
rect 38 103 67 109
rect 117 128 146 139
rect 117 111 123 128
rect 142 111 146 128
rect 117 103 146 111
rect 35 64 67 70
rect 35 47 42 64
rect 60 47 67 64
rect 35 34 67 47
rect 117 34 139 70
rect 189 64 223 70
rect 189 47 196 64
rect 216 47 223 64
rect 189 34 223 47
<< mvpdiffc >>
rect 42 109 60 126
rect 123 111 142 128
rect 42 47 60 64
rect 196 47 216 64
<< mvnsubdiff >>
rect 189 128 223 142
rect 189 110 196 128
rect 216 110 223 128
rect 189 98 223 110
<< mvnsubdiffcont >>
rect 196 110 216 128
<< poly >>
rect 67 139 117 152
rect 67 95 117 103
rect 0 78 117 95
rect 154 86 173 164
rect 67 70 117 78
rect 139 70 189 86
rect 67 21 117 34
rect 139 1 189 34
<< locali >>
rect 123 128 143 136
rect 34 109 42 126
rect 60 109 68 126
rect 142 111 143 128
rect 123 97 143 111
rect 123 80 124 97
rect 141 80 143 97
rect 123 76 143 80
rect 195 128 217 136
rect 195 110 196 128
rect 216 110 217 128
rect 195 94 217 110
rect 195 77 197 94
rect 214 77 217 94
rect 196 74 217 77
rect 196 64 216 74
rect 34 47 42 64
rect 60 47 68 64
rect 196 39 216 47
<< viali >>
rect 124 80 141 97
rect 197 77 214 94
<< metal1 >>
rect 123 105 139 191
rect 163 117 179 191
rect 204 140 220 191
rect 204 131 221 140
rect 162 105 179 117
rect 123 100 144 105
rect 121 97 144 100
rect 121 80 124 97
rect 141 80 144 97
rect 121 76 144 80
rect 123 74 143 76
rect 123 1 139 74
rect 160 6 179 105
rect 193 126 221 131
rect 193 94 220 126
rect 193 77 197 94
rect 214 77 220 94
rect 193 71 220 77
rect 204 1 220 71
<< metal2 >>
rect 0 99 9 117
rect 39 99 256 117
rect 38 56 256 74
use sky130_hilas_li2m2  sky130_hilas_li2m2_0
timestamp 1634057699
transform 1 0 23 0 -1 60
box 0 0 34 33
use sky130_hilas_li2m2  sky130_hilas_li2m2_1
timestamp 1634057699
transform 1 0 23 0 -1 115
box 0 0 34 33
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
