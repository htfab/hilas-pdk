VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
  WIDTH 0.030000 ;
  SPACING 0.040000 ;
  DIRECTION HORIZONTAL ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  SPACING 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  SPACING 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  SPACING 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  SPACING 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO sky130_hilas_pfetdevice01a
  CLASS BLOCK ;
  FOREIGN sky130_hilas_pfetdevice01a ;
  ORIGIN 0.800 0.420 ;
  SIZE 1.610 BY 0.850 ;
  OBS
      LAYER nwell ;
        RECT -0.800 -0.420 0.810 0.430 ;
  END
END sky130_hilas_pfetdevice01a
END LIBRARY

