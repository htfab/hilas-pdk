magic
tech sky130A
timestamp 1628178864
<< error_p >>
rect -465 248 -463 298
rect -423 248 -421 298
rect -330 248 -327 298
rect -288 248 -285 298
rect -465 169 -463 219
rect -423 169 -421 219
rect -330 169 -327 219
rect -288 169 -285 219
rect -463 142 -423 144
rect -327 142 -288 144
rect -256 142 -249 144
rect -222 111 -172 117
rect -150 111 -100 117
rect -222 69 -172 75
rect -150 69 -100 75
<< nwell >>
rect -364 42 -33 359
<< mvnmos >>
rect -463 248 -423 298
rect -463 169 -423 219
<< mvpmos >>
rect -327 248 -288 298
rect -327 169 -288 219
rect -224 142 -173 326
rect -222 75 -172 111
rect -150 75 -100 111
<< mvndiff >>
rect -463 321 -423 326
rect -463 304 -452 321
rect -434 304 -423 321
rect -463 298 -423 304
rect -463 242 -423 248
rect -463 225 -453 242
rect -434 225 -423 242
rect -463 219 -423 225
rect -463 163 -423 169
rect -463 146 -452 163
rect -434 146 -423 163
rect -463 142 -423 146
<< mvpdiff >>
rect -327 321 -288 326
rect -327 304 -316 321
rect -299 304 -288 321
rect -327 298 -288 304
rect -256 305 -224 326
rect -256 288 -249 305
rect -232 288 -224 305
rect -256 271 -224 288
rect -256 254 -249 271
rect -232 254 -224 271
rect -327 242 -288 248
rect -327 225 -316 242
rect -299 225 -288 242
rect -327 219 -288 225
rect -256 237 -224 254
rect -256 220 -249 237
rect -232 220 -224 237
rect -256 203 -224 220
rect -256 186 -249 203
rect -232 186 -224 203
rect -256 169 -224 186
rect -327 163 -288 169
rect -327 146 -316 163
rect -299 146 -288 163
rect -327 142 -288 146
rect -256 152 -249 169
rect -232 152 -224 169
rect -256 142 -224 152
rect -173 304 -145 326
rect -173 287 -166 304
rect -149 287 -145 304
rect -173 270 -145 287
rect -173 253 -166 270
rect -149 253 -145 270
rect -173 236 -145 253
rect -173 219 -166 236
rect -149 219 -145 236
rect -173 202 -145 219
rect -173 185 -166 202
rect -149 185 -145 202
rect -173 168 -145 185
rect -173 151 -166 168
rect -149 151 -145 168
rect -173 142 -145 151
rect -256 105 -222 111
rect -256 88 -247 105
rect -229 88 -222 105
rect -256 75 -222 88
rect -172 75 -150 111
rect -100 105 -66 111
rect -100 88 -93 105
rect -73 88 -66 105
rect -100 75 -66 88
<< mvndiffc >>
rect -452 304 -434 321
rect -453 225 -434 242
rect -452 146 -434 163
<< mvpdiffc >>
rect -316 304 -299 321
rect -249 288 -232 305
rect -249 254 -232 271
rect -316 225 -299 242
rect -249 220 -232 237
rect -249 186 -232 203
rect -316 146 -299 163
rect -249 152 -232 169
rect -166 287 -149 304
rect -166 253 -149 270
rect -166 219 -149 236
rect -166 185 -149 202
rect -166 151 -149 168
rect -247 88 -229 105
rect -93 88 -73 105
<< mvnsubdiff >>
rect -100 169 -66 183
rect -100 151 -93 169
rect -73 151 -66 169
rect -100 139 -66 151
<< mvnsubdiffcont >>
rect -93 151 -73 169
<< poly >>
rect -224 326 -173 339
rect -476 248 -463 298
rect -423 248 -327 298
rect -288 248 -275 298
rect -476 169 -463 219
rect -423 169 -327 219
rect -288 169 -275 219
rect -133 248 -98 256
rect -133 231 -121 248
rect -104 231 -98 248
rect -133 223 -98 231
rect -133 222 -104 223
rect -133 193 -106 222
rect -476 134 -257 136
rect -224 134 -173 142
rect -476 119 -172 134
rect -129 127 -106 193
rect -129 125 -100 127
rect -222 111 -172 119
rect -150 111 -100 125
rect -222 60 -172 75
rect -150 60 -100 75
<< polycont >>
rect -121 231 -104 248
<< locali >>
rect -460 304 -452 321
rect -434 304 -426 321
rect -324 304 -316 321
rect -299 304 -291 321
rect -249 305 -232 313
rect -249 271 -232 288
rect -461 225 -453 242
rect -434 225 -426 242
rect -324 225 -316 242
rect -299 225 -291 242
rect -249 237 -232 254
rect -249 203 -232 220
rect -249 169 -232 186
rect -461 146 -452 163
rect -434 146 -426 163
rect -324 146 -316 163
rect -299 146 -291 163
rect -249 144 -232 152
rect -166 270 -149 287
rect -166 236 -149 253
rect -130 248 -103 256
rect -130 231 -121 248
rect -104 231 -103 248
rect -130 223 -103 231
rect -166 202 -149 219
rect -129 219 -109 223
rect -129 200 -128 219
rect -110 200 -109 219
rect -129 194 -109 200
rect -129 193 -110 194
rect -166 168 -149 185
rect -93 176 -72 177
rect -166 143 -149 151
rect -94 169 -72 176
rect -94 151 -93 169
rect -73 151 -72 169
rect -94 135 -72 151
rect -94 118 -92 135
rect -75 118 -72 135
rect -93 115 -72 118
rect -93 105 -73 115
rect -256 88 -247 105
rect -229 88 -221 105
rect -93 80 -73 88
<< viali >>
rect -166 304 -148 323
rect -128 200 -110 219
rect -92 118 -75 135
rect -274 88 -256 105
<< metal1 >>
rect -169 323 -145 329
rect -169 304 -166 323
rect -148 304 -145 323
rect -169 291 -145 304
rect -126 248 -110 350
rect -130 224 -107 248
rect -130 223 -106 224
rect -131 219 -106 223
rect -131 200 -128 219
rect -110 200 -106 219
rect -131 196 -106 200
rect -129 193 -107 196
rect -281 126 -250 129
rect -281 100 -278 126
rect -252 100 -250 126
rect -281 88 -274 100
rect -256 88 -250 100
rect -281 85 -250 88
rect -129 48 -110 193
rect -85 181 -69 350
rect -85 172 -68 181
rect -96 167 -68 172
rect -96 135 -69 167
rect -96 118 -92 135
rect -75 118 -69 135
rect -96 112 -69 118
rect -85 48 -69 112
<< via1 >>
rect -278 105 -252 126
rect -278 100 -274 105
rect -274 100 -256 105
rect -256 100 -252 105
<< metal2 >>
rect -281 126 -250 129
rect -281 100 -278 126
rect -252 115 -250 126
rect -252 100 -33 115
rect -281 97 -33 100
rect -281 96 -250 97
<< end >>
