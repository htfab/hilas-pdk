magic
tech sky130A
timestamp 1607392100
<< error_s >>
rect -91 192 -62 210
rect 155 190 184 206
rect 234 190 263 206
rect 313 190 342 206
rect 392 190 421 206
rect -91 160 -90 161
rect -63 160 -62 161
rect -141 131 -123 160
rect -92 159 -61 160
rect -91 150 -62 159
rect -91 141 -81 150
rect -72 141 -62 150
rect -91 132 -62 141
rect -92 131 -61 132
rect -30 131 -12 160
rect 155 156 156 157
rect 183 156 184 157
rect 234 156 235 157
rect 262 156 263 157
rect 313 156 314 157
rect 341 156 342 157
rect 392 156 393 157
rect 420 156 421 157
rect -91 130 -90 131
rect -63 130 -62 131
rect 105 127 123 156
rect 154 155 185 156
rect 233 155 264 156
rect 312 155 343 156
rect 391 155 422 156
rect 155 148 184 155
rect 234 148 263 155
rect 313 148 342 155
rect 392 148 421 155
rect 155 134 165 148
rect 412 134 421 148
rect 155 128 184 134
rect 234 128 263 134
rect 313 128 342 134
rect 392 128 421 134
rect 154 127 185 128
rect 233 127 264 128
rect 312 127 343 128
rect 391 127 422 128
rect 454 127 471 156
rect 488 134 490 135
rect 155 126 156 127
rect 183 126 184 127
rect 234 126 235 127
rect 262 126 263 127
rect 313 126 314 127
rect 341 126 342 127
rect 392 126 393 127
rect 420 126 421 127
rect -91 81 -62 99
rect 155 77 184 92
rect 234 77 263 92
rect 313 77 342 92
rect 392 77 421 92
rect -91 40 -62 58
rect 155 43 184 59
rect 234 43 263 59
rect 313 43 342 59
rect 392 43 421 59
rect 155 9 156 10
rect 183 9 184 10
rect 234 9 235 10
rect 262 9 263 10
rect 313 9 314 10
rect 341 9 342 10
rect 392 9 393 10
rect 420 9 421 10
rect -91 8 -90 9
rect -63 8 -62 9
rect -141 -21 -123 8
rect -92 7 -61 8
rect -91 -2 -62 7
rect -91 -11 -81 -2
rect -72 -11 -62 -2
rect -91 -20 -62 -11
rect -92 -21 -61 -20
rect -30 -21 -12 8
rect 105 -20 123 9
rect 154 8 185 9
rect 233 8 264 9
rect 312 8 343 9
rect 391 8 422 9
rect 155 1 184 8
rect 234 1 263 8
rect 313 1 342 8
rect 392 1 421 8
rect 155 -13 165 1
rect 412 -13 421 1
rect 155 -19 184 -13
rect 234 -19 263 -13
rect 313 -19 342 -13
rect 392 -19 421 -13
rect 154 -20 185 -19
rect 233 -20 264 -19
rect 312 -20 343 -19
rect 391 -20 422 -19
rect 454 -20 471 9
rect 483 -17 496 -13
rect 497 -17 510 -12
rect 483 -20 510 -17
rect 155 -21 156 -20
rect 183 -21 184 -20
rect 234 -21 235 -20
rect 262 -21 263 -20
rect 313 -21 314 -20
rect 341 -21 342 -20
rect 392 -21 393 -20
rect 420 -21 421 -20
rect -91 -22 -90 -21
rect -63 -22 -62 -21
rect -91 -71 -62 -53
rect 155 -70 184 -55
rect 234 -70 263 -55
rect 313 -70 342 -55
rect 392 -70 421 -55
rect -91 -105 -62 -87
rect 155 -104 184 -88
rect 234 -104 263 -88
rect 313 -104 342 -88
rect 392 -104 421 -88
rect -91 -137 -90 -136
rect -63 -137 -62 -136
rect -141 -166 -123 -137
rect -92 -138 -61 -137
rect -91 -147 -62 -138
rect -91 -156 -81 -147
rect -72 -156 -62 -147
rect -91 -165 -62 -156
rect -92 -166 -61 -165
rect -30 -166 -12 -137
rect 155 -138 156 -137
rect 183 -138 184 -137
rect 234 -138 235 -137
rect 262 -138 263 -137
rect 313 -138 314 -137
rect 341 -138 342 -137
rect 392 -138 393 -137
rect 420 -138 421 -137
rect -91 -167 -90 -166
rect -63 -167 -62 -166
rect 105 -167 123 -138
rect 154 -139 185 -138
rect 233 -139 264 -138
rect 312 -139 343 -138
rect 391 -139 422 -138
rect 155 -146 184 -139
rect 234 -146 263 -139
rect 313 -146 342 -139
rect 392 -146 421 -139
rect 155 -160 165 -146
rect 412 -160 421 -146
rect 155 -166 184 -160
rect 234 -166 263 -160
rect 313 -166 342 -160
rect 392 -166 421 -160
rect 154 -167 185 -166
rect 233 -167 264 -166
rect 312 -167 343 -166
rect 391 -167 422 -166
rect 454 -167 471 -138
rect 155 -168 156 -167
rect 183 -168 184 -167
rect 234 -168 235 -167
rect 262 -168 263 -167
rect 313 -168 314 -167
rect 341 -168 342 -167
rect 392 -168 393 -167
rect 420 -168 421 -167
rect -91 -216 -62 -198
rect 155 -217 184 -202
rect 234 -217 263 -202
rect 313 -217 342 -202
rect 392 -217 421 -202
rect -91 -259 -62 -241
rect 155 -251 184 -235
rect 234 -251 263 -235
rect 313 -251 342 -235
rect 392 -251 421 -235
rect 155 -285 156 -284
rect 183 -285 184 -284
rect 234 -285 235 -284
rect 262 -285 263 -284
rect 313 -285 314 -284
rect 341 -285 342 -284
rect 392 -285 393 -284
rect 420 -285 421 -284
rect -91 -291 -90 -290
rect -63 -291 -62 -290
rect -141 -320 -123 -291
rect -92 -292 -61 -291
rect -91 -301 -62 -292
rect -91 -310 -81 -301
rect -72 -310 -62 -301
rect -91 -319 -62 -310
rect -92 -320 -61 -319
rect -30 -320 -12 -291
rect 105 -314 123 -285
rect 154 -286 185 -285
rect 233 -286 264 -285
rect 312 -286 343 -285
rect 391 -286 422 -285
rect 155 -293 184 -286
rect 234 -293 263 -286
rect 313 -293 342 -286
rect 392 -293 421 -286
rect 155 -307 165 -293
rect 412 -307 421 -293
rect 155 -313 184 -307
rect 234 -313 263 -307
rect 313 -313 342 -307
rect 392 -313 421 -307
rect 154 -314 185 -313
rect 233 -314 264 -313
rect 312 -314 343 -313
rect 391 -314 422 -313
rect 454 -314 471 -285
rect 155 -315 156 -314
rect 183 -315 184 -314
rect 234 -315 235 -314
rect 262 -315 263 -314
rect 313 -315 314 -314
rect 341 -315 342 -314
rect 392 -315 393 -314
rect 420 -315 421 -314
rect -91 -321 -90 -320
rect -63 -321 -62 -320
rect -91 -370 -62 -352
rect 155 -364 184 -349
rect 234 -364 263 -349
rect 313 -364 342 -349
rect 392 -364 421 -349
<< nwell >>
rect 632 -72 667 -71
rect 632 -88 649 -72
rect 666 -88 667 -72
<< poly >>
rect 469 147 489 151
rect -19 114 130 138
rect 469 135 488 147
rect -19 5 128 29
rect 469 -9 488 8
rect 649 -72 667 -71
rect 665 -88 667 -72
rect -19 -175 130 -151
rect 469 -167 488 -150
rect -19 -295 132 -271
rect 469 -309 488 -292
<< polycont >>
rect 632 -88 649 -71
<< locali >>
rect 623 -88 632 -71
<< viali >>
rect 649 -88 667 -71
<< metal1 >>
rect -90 -382 -63 223
rect 654 -68 667 -66
rect 646 -71 670 -68
rect 646 -88 649 -71
rect 667 -88 670 -71
rect 646 -91 670 -88
rect 656 -95 667 -91
<< metal2 >>
rect -191 166 497 173
rect -191 155 500 166
rect -191 112 710 130
rect -191 24 497 30
rect -191 12 500 24
rect -191 -20 496 -13
rect -191 -31 500 -20
rect -191 -146 500 -129
rect -191 -188 500 -171
rect -191 -286 500 -269
rect -191 -330 500 -313
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_3
timestamp 1607262215
transform 1 0 -79 0 1 -327
box -62 -43 67 86
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_2
timestamp 1607262215
transform 1 0 -79 0 1 -173
box -62 -43 67 86
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_3
timestamp 1607261501
transform 1 0 609 0 1 -328
box -521 -54 -121 110
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_2
timestamp 1607261501
transform 1 0 609 0 1 -181
box -521 -54 -121 110
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_1
timestamp 1607386385
transform 1 0 777 0 1 -428
box -289 47 -33 232
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_2
timestamp 1607386385
transform 1 0 777 0 -1 -31
box -289 47 -33 232
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_1
timestamp 1607262215
transform 1 0 -79 0 1 -28
box -62 -43 67 86
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_1
timestamp 1607261501
transform 1 0 609 0 1 -34
box -521 -54 -121 110
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_0
timestamp 1607386385
transform 1 0 777 0 1 -128
box -289 47 -33 232
use sky130_hilas_nOverlapCap01  sky130_hilas_nOverlapCap01_0
timestamp 1607262215
transform 1 0 -79 0 1 124
box -62 -43 67 86
use sky130_hilas_overlapCap02a  sky130_hilas_overlapCap02a_0
timestamp 1607261501
transform 1 0 609 0 1 113
box -521 -54 -121 110
use sky130_hilas_horizPcell01  sky130_hilas_horizPcell01_3
timestamp 1607386385
transform 1 0 777 0 -1 270
box -289 47 -33 232
<< end >>
